module poseONE_tb;
	reg clock;
	reg validIn;
	reg reset;
	reg signed [12:0] Rx, Ry;
	wire [15:0] LUTin;
	wire signed [12:0] atan;
	wire validOut;

 	localparam [17:0]
	bx1 = 18'b11011110_1000000000, by1 = 18'b01001001_0000000000, bz1 = 18'b00000000_0000000000,
 	bx2 = 18'b00100001_1000000000, by2 = 18'b01001001_0000000000, bz2 = 18'b00000000_0000000000,
 	bx3 = 18'b01010000_0000000000, by3 = 18'b11111000_1000000000, bz3 = 18'b00000000_0000000000,
 	bx4 = 18'b00101110_1000000000, by4 = 18'b10111110_1000000000, bz4 = 18'b00000000_0000000000,
 	bx5 = 18'b11010001_1000000000, by5 = 18'b10111110_1000000000, bz5 = 18'b00000000_0000000000,
 	bx6 = 18'b10110000_0000000000, by6 = 18'b11111000_1000000000, bz6 = 18'b00000000_0000000000,
 	px1 = 18'b11010100_1110011001, py1 = 18'b00100111_0100110011, pz1 = 18'b00000000_0000000000,
 	px2 = 18'b00101011_0001100110, py2 = 18'b00100111_0100110011, pz2 = 18'b00000000_0000000000,
 	px3 = 18'b00110111_1001100110, py3 = 18'b00010001_1011001100, pz3 = 18'b00000000_0000000000,
 	px4 = 18'b00001100_1000000000, py4 = 18'b11000111_0000000000, pz4 = 18'b00000000_0000000000,
 	px5 = 18'b11110011_1000000000, py5 = 18'b11000111_0000000000, pz5 = 18'b00000000_0000000000,
	px6 = 18'b11001000_0110011001, py6 = 18'b00010001_1011001100, pz6 = 18'b00000000_0000000000;

	localparam [12:0] 
	ZERO = 13'b000_0000000000, 
	THIRTY = 13'b000_0010101010,
	NTHIRTY = 13'b111_1101010101;

	// BETAS = 90 90 330 330 210 210
	poseONE #(.BETA(90)) 
		uut(.clock(clock),
			.validIn(validIn),
			.reset(reset),
			.bx(bx1),.by(by1),.bz(bz1),
			.px(px1),.py(py1),.pz(pz1),
			.Rx(Rx),.Ry(Ry),
			.LUTin(LUTin),
			.atan(atan),
			.validOut(validOut));

	always #5 clock <= ~clock;

    initial begin
        clock = 0;
        validIn = 0;
        reset = 0;
        Rx = ZERO;
        Ry = ZERO;
        #100
        reset = 1;
        #10
        reset = 0;
        Rx = NTHIRTY; // -30 degrees
        Ry = THIRTY; // 30 degrees
        #5
        validIn = 1;
        #5
        validIn = 0;
    end

endmodule
