`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/08/2018 11:35:18 PM
// Design Name: 
// Module Name: dp_3x1_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module dp_3x1_tb;

    parameter A_WIDTH = 18;
    parameter B_WIDTH = 18;

    reg clock;
    reg validIn;
    reg reset;
    reg [A_WIDTH-1:0] A1, A2, A3;
    reg [B_WIDTH-1:0] B1, B2, B3;
    wire [A_WIDTH + B_WIDTH:0] dp;
    wire validOut;

    localparam [17:0]
    bx1 = 18'b11011110_1000000000, by1 = 18'b01001001_0000000000, bz1 = 18'b00000000_0000000000,
    bx2 = 18'b00100001_1000000000, by2 = 18'b01001001_0000000000, bz2 = 18'b00000000_0000000000,
    bx3 = 18'b01010000_0000000000, by3 = 18'b11111000_1000000000, bz3 = 18'b00000000_0000000000,
    bx4 = 18'b00101110_1000000000, by4 = 18'b10111110_1000000000, bz4 = 18'b00000000_0000000000,
    bx5 = 18'b11010001_1000000000, by5 = 18'b10111110_1000000000, bz5 = 18'b00000000_0000000000,
    bx6 = 18'b10110000_0000000000, by6 = 18'b11111000_1000000000, bz6 = 18'b00000000_0000000000,
    px1 = 18'b11010100_1110011001, py1 = 18'b00100111_0100110011, pz1 = 18'b00000000_0000000000,
    px2 = 18'b00101011_0001100110, py2 = 18'b00100111_0100110011, pz2 = 18'b00000000_0000000000,
    px3 = 18'b00110111_1001100110, py3 = 18'b00010001_1011001100, pz3 = 18'b00000000_0000000000,
    px4 = 18'b00001100_1000000000, py4 = 18'b11000111_0000000000, pz4 = 18'b00000000_0000000000,
    px5 = 18'b11110011_1000000000, py5 = 18'b11000111_0000000000, pz5 = 18'b00000000_0000000000,
    px6 = 18'b11001000_0110011001, py6 = 18'b00010001_1011001100, pz6 = 18'b00000000_0000000000;

    localparam [15:0] // Computing using Rx = -30deg and Ry = 30deg
    R11 = 16'b00_11011101111110, R12 = 16'b11_11101110111000, R13 = 16'b00_00111111110000,
    R21 = 16'b00_00000000000000, R22 = 16'b00_11011101100101, R23 = 16'b00_10000000001110,
    R31 = 16'b11_10000000011101, R32 = 16'b11_10111111110111, R33 = 16'b00_11101110111000;
    
    dp_3x1 #(.A_WIDTH(A_WIDTH), .B_WIDTH(B_WIDTH))
        uut(.clock(clock),
            .validIn(validIn),
            .reset(reset),
            .A1(A1),
            .A2(A2),
            .A3(A3),
            .B1(B1),
            .B2(B2),
            .B3(B3),
            .dp(dp),
            .validOut(validOut));
    
    always #5 clock <= ~clock;
    
    initial begin
        clock = 0;
        validIn = 0;
        reset = 0;
        #100
        reset = 1;
        #10
        reset = 0;
        A1 = R11 << 2;
        A2 = R12 << 2;
        A3 = R13 << 2;
        B1 = px1;
        B2 = px2;
        B3 = px3;
        #5
        validIn = 1;
        #5
        validIn = 0;
    end
        
endmodule
